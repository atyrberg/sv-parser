module mod_w_inc ();
    // Including on line 3
    `include "test3.svh"
    logic not_in_inc_file = 2;
endmodule
