// Line 1
localparam INC_FILE = 1;
// Line 3
